library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all; -- BIBLIOTECA PADRÃO

entity banco_registradores is
	Port (	i_CLK  	: in std_logic;
    		i_RSTn	: in std_logic;
            i_WRena	: in std_logic;
            i_WRaddr: in std_logic_vector(4 downto 0);
    		i_RS1 	: in std_logic_vector(4 downto 0);
            i_RS2 	: in std_logic_vector(4 downto 0);
            i_DATA 	: in std_logic_vector(31 downto 0);
            o_RS1 	: out std_logic_vector(31 downto 0);
            o_RS2 	: out std_logic_vector(31 downto 0)
         );
end banco_registradores;

architecture arch_1 of banco_registradores is
	type t_MEMORIA is array(0 to 31) of std_logic_vector(31 downto 0);
    signal w_REG : t_MEMORIA := (others => (others => '0'));

begin
    process( i_CLK, i_RSTn )
    begin
        if i_RSTn = '0' then
            w_REG <= (others => (others => '0'));
        elsif rising_edge(i_CLK) then               
            if i_WRena = '1' and i_WRaddr /= "00000" then
                -- CONVERSÃO EXPLÍCITA E SEGURA
                w_REG(to_integer(unsigned(i_WRaddr))) <= i_DATA;
            end if;
        end if;
    end process;

    -- Leituras combinacionais (assíncronas)
    o_RS1 <= w_REG(to_integer(unsigned(i_RS1))) when i_RS1 /= "00000" else (others => '0');
    o_RS2 <= w_REG(to_integer(unsigned(i_RS2))) when i_RS2 /= "00000" else (others => '0');

end arch_1;
